Ring Oscillator Design

.SUBCKT INVERTER  INPUT OUTPUT
.ENDS INVERTER