Ring Oscillator Design

.SUBCKT INVERTER IN OUT VDD DGND ;
.include cmosedu_models.txt
M1 OUT IN VDD  VDD  P_50n    ;M1 OUT IN VDD  VDD  MOSP
M2 OUT IN DGND DGND N_50n    ;M2 OUT IN DGND DGND MOSN
.ENDS INVERTER

X01 IN01 IN02 VDD DGND INVERTER
X02 IN02 IN03 VDD DGND INVERTER
X03 IN03 IN04 VDD DGND INVERTER
X04 IN04 IN05 VDD DGND INVERTER
X05 IN05 IN06 VDD DGND INVERTER
X06 IN06 IN07 VDD DGND INVERTER
X07 IN07 IN08 VDD DGND INVERTER
X08 IN08 IN09 VDD DGND INVERTER
X09 IN09 IN10 VDD DGND INVERTER
X10 IN10 IN11 VDD DGND INVERTER
X11 IN11 IN12 VDD DGND INVERTER
X12 IN12 IN13 VDD DGND INVERTER
X13 IN13 IN14 VDD DGND INVERTER
X14 IN14 IN15 VDD DGND INVERTER
X15 IN15 IN16 VDD DGND INVERTER
X16 IN16 IN17 VDD DGND INVERTER
X17 IN17 IN01 VDD DGND INVERTER

.control
echo ******************************************
echo *** Ring Oscillator Simulation Started ***
echo ******************************************
run
echo *******************************************
echo *** Ring Oscillator Simulation Finished ***
echo *******************************************
.endc
.END         ; End of the file