Ring Oscillator Design

.SUBCKT INVERTER IN OUT VDD DGND
M1 OUT IN VDD  VDD  MOSP
M2 OUT IN DGND DGND MOSN
.ENDS INVERTER

.END         ; End of the file