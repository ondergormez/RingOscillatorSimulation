Ring Oscillator Design


VDD NVDD GND DC 5

.SUBCKT INVERTER IN OUT VDD DGND                                                ;Inverter Sub circuit
.include cmosedu_models.txt
M1 OUT IN VDD  VDD  P_50n    ;M1 OUT IN VDD  VDD  MOSP
M2 OUT IN DGND DGND N_50n    ;M2 OUT IN DGND DGND MOSN
.ENDS INVERTER

X01 IN01 IN02 NVDD GND INVERTER                                                ;TODO: Change NVDD to VDD and observe the simulation result!
X02 IN02 IN03 NVDD GND INVERTER
X03 IN03 IN04 NVDD GND INVERTER
X04 IN04 IN05 NVDD GND INVERTER
X05 IN05 IN06 NVDD GND INVERTER
X06 IN06 IN07 NVDD GND INVERTER
X07 IN07 IN08 NVDD GND INVERTER
X08 IN08 IN09 NVDD GND INVERTER
X09 IN09 IN10 NVDD GND INVERTER
X10 IN10 IN11 NVDD GND INVERTER
X11 IN11 IN12 NVDD GND INVERTER
X12 IN12 IN13 NVDD GND INVERTER
X13 IN13 IN14 NVDD GND INVERTER
X14 IN14 IN15 NVDD GND INVERTER
X15 IN15 IN16 NVDD GND INVERTER
X16 IN16 IN17 NVDD GND INVERTER
X17 IN17 IN01 NVDD GND INVERTER

.control
echo ******************************************
echo *** Ring Oscillator Simulation Started ***
echo ******************************************
run
echo *******************************************
echo *** Ring Oscillator Simulation Finished ***
echo *******************************************
.endc
.END         ; End of the file